entity hallo is 
end hallo;

architecture sim of hallo is
 begin

  process
  begin
    report "i hallo venkatesh";
  end process;

 
end sim;
